interface comparator_if(input logic clk, reset);
  logic ip1, ip2;
  logic gt,eq,lt;
  
  /*clocking driver_cb @(posedge clk);
    default input #1 output #1;
  endclocking
  */
endinterface
